`timescale 1ps / 1ps
module tb_syn_ksa();

// Your testbench goes here.

endmodule: tb_syn_ksa
